II* 
             �       
     .       *      II* 
   
* 
I  3I*